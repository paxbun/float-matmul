// Copyright (c) 2021 Chanjung Kim (paxbun). All rights reserved.
// Licensed under the MIT License.

`ifndef LZC_MACROS_VH
`define LZC_MACROS_VH

`define LZC_PARAMS              \
    parameter INPUT_WIDTH = 26, \
    parameter OUTPUT_WIDTH = 5, \
    parameter OUTPUT_STEP = 1,  \
    parameter OUTPUT_BIAS = 0

`endif